always @(*) begin
   case (function)
      0:
        default:
